VIEW   1, 1, 0, 0, 0, 1, 0, 0, 0, 1
VIEW   2, 1, 0, 0, 0, 0, -1, 0, 1, 0
VIEW   3, -1, 0, 0, 0, 0, 1, 0, 1, 0
VIEW   4, -1, 0, 0, 0, 1, 0, 0, 0, -1
VIEW   5, 0, 0, 1, 1, 0, 0, 0, 1, 0
VIEW   6, 0, 0, -1, -1, 0, 0, 0, 1, 0
VIEW   7, 0.7071068, -0.4082483, 0.5773503, 0.7071068, 0.4082483, -0.5773503, 0, 0.8164966, 0.5773503
VIEW   8, 0.5, 0.5, 0.707107, -0.853553, 0.146447, 0.5, 0.146447, -0.853553, 0.5
VIEW   9, 1, 0, 0, 0, -1, 0, 0, 0, -1
VIEW   10, 0.8660254, 0, -0.5, -0.5, 0, -0.8660254, 0, 1, 0
VIEW   11, 0.5, 0, 0.8660254, 0.8660254, 0, -0.5, 0, 1, 0
VIEW   12, 0.8660254, 0, 0.5, 0.5, 0, -0.8660254, 0, 1, 0
LINE   2.133975, 0, 18.75, 3, 0, 18.25, 11, 101, 1
LINE   3.464102, 2, 9, 8.660254, 5, 13, 12, 43, 1
LINE   0.01, 12, 9, 0.01, -12, 9, 4, 41, 1
LINE   15, -12, 9, 0.01, -12, 9, 4, 41, 1
LINE   10, 0, 13, 10, 0, 15, 12, 43, 1
LINE   10, 0, 15, 4, 2.220446E-016, 19, 12, 43, 1
LINE   15, -12, 9, 15, 24.90126, 9, 4, 41, 1
LINE   4, 0, 9, 10, 0, 13, 12, 43, 1
LINE   4, 0, 9, 0, 0, 9, 12, 43, 1
LINE   4, 0, 19, 0, 0, 19, 12, 43, 1
CIRCLE -13, 14, 12, 2.99, 2, 12, 36, 1
CIRCLE -17.5, -9, 9, 1.5, 1, 12, 36, 1
CIRCLE 0, 14, -20, 1, 5, 12, 36, 1
CIRCLE -9, 17.5, -12, 1, 2, 12, 36, 1
CIRCLE -17.5, 9, 9, 1.5, 1, 12, 36, 1
LINE   -0.01, -12, 9, -20, -12, 9, 9, 36, 1
LINE   -0.01, 12, 9, -0.01, -12, 9, 9, 36, 1
LINE   -20, 12, 9, -0.01, 12, 9, 9, 36, 1
LINE   -20, -12, 9, -20, 12, 9, 9, 36, 1
LINE   0, 0, 19, 0, 0, 9, 12, 43, 1
LINE   3.332996, 1.924306, 19, 2.223076, 1.283494, 19, 11, 101, 1
ARC    3.848612, 18.5, 2.220446E-016, 0.5, 56.30993, 90, 12, 10, 101, 1
LINE   3.573188, 2.062981, 18.91603, 8.467434, 4.888675, 15.14843, 10, 101, 1
ARC    9.5, 14.73241, 0, 0.5, 0, 56.30993, 12, 10, 101, 1
LINE   8.660254, 5, 14.73241, 8.660254, 5, 13.26759, 10, 101, 1
ARC    9.5, 13.26759, 0, 0.5, 303.6901, 360, 12, 10, 101, 1
LINE   8.467434, 4.888675, 12.85157, 3.573188, 2.062981, 9.083975, 10, 101, 1
ARC    3.848612, 9.5, 0, 0.5, 270, 303.6901, 12, 10, 101, 1
LINE   2.223076, 1.283494, 9, 3.332996, 1.924306, 9, 11, 101, 1
LINE   2.598076, 1.5, 9.25, 2.223076, 1.283494, 9, 11, 101, 1
LINE   1.848076, 1.066987, 9.75, 2.598076, 1.5, 9.25, 11, 101, 1
LINE   2.598076, 1.5, 10.25, 1.848076, 1.066987, 9.75, 11, 101, 1
LINE   2.598076, 1.5, 10.25, 1.848076, 1.066987, 10.75, 11, 101, 1
LINE   2.598076, 1.5, 11.25, 1.848076, 1.066987, 10.75, 11, 101, 1
LINE   1.848076, 1.066987, 11.75, 2.598076, 1.5, 11.25, 11, 101, 1
LINE   2.598076, 1.5, 12.25, 1.848076, 1.066987, 11.75, 11, 101, 1
LINE   1.848076, 1.066987, 12.75, 2.598076, 1.5, 12.25, 11, 101, 1
LINE   2.598076, 1.5, 13.25, 1.848076, 1.066987, 12.75, 11, 101, 1
LINE   1.848076, 1.066987, 13.75, 2.598076, 1.5, 13.25, 11, 101, 1
LINE   2.598076, 1.5, 14.25, 1.848076, 1.066987, 13.75, 11, 101, 1
LINE   1.848076, 1.066987, 14.75, 2.598076, 1.5, 14.25, 11, 101, 1
LINE   2.598076, 1.5, 15.25, 1.848076, 1.066987, 14.75, 11, 101, 1
LINE   1.848076, 1.066987, 15.75, 2.598076, 1.5, 15.25, 11, 101, 1
LINE   2.598076, 1.5, 16.25, 1.848076, 1.066987, 15.75, 11, 101, 1
LINE   2.598076, 1.5, 16.25, 1.848076, 1.066987, 16.75, 11, 101, 1
LINE   2.598076, 1.5, 17.25, 1.848076, 1.066987, 16.75, 11, 101, 1
LINE   1.848076, 1.066987, 17.75, 2.598076, 1.5, 17.25, 11, 101, 1
LINE   2.598076, 1.5, 18.25, 1.848076, 1.066987, 17.75, 11, 101, 1
LINE   1.848076, 1.066987, 18.75, 2.598076, 1.5, 18.25, 11, 101, 1
LINE   2.223076, 1.283494, 19, 1.848076, 1.066987, 18.75, 11, 101, 1
CIRCLE 11.5, 24.90126, 9, 1.5, 1, 14, 41, 1
LINE   0.01, 12, 9, 8.468911, 26.65126, 9, 4, 102, 1
ARC    11.5, 24.90126, 9, 3.5, 0, 150, 1, 4, 102, 1
CIRCLE 5.5, 14.50896, 9, 1.5, 1, 14, 41, 1
LINE   0.7032248, 14.2007, 14, 8.035898, 26.90126, 14, 10, 43, 1
LINE   0.7032248, 14.2007, 14, 15.5, 7.300852, 14, 10, 43, 1
LINE   15.5, 24.90126, 14, 15.5, 7.300852, 14, 4, 102, 1
ARC    11.5, 24.90126, 14, 4, 360, 510, 1, 10, 43, 1
